Unity-gain feedback op-amp

* Circuit Description
* We will used voltage control current source and voltage control voltage source
* to make a small signal model

* Add the subcircuit
.LIB Non_ideal_op_amp.lib

* Subcircuit Inantiation
Xop_amp 1 2 1 small_signal_opamp

* parametric sweep for RF
*.STEP PARAM RFED LIST 4k, 9k
* Signal sources
*2 Vin 2 0 DC 1
*3-6Vsig 2 0 SIN(0 1 {freq} 0 0 0)
Vin 2 0 AC 1
* Circuit elements
* R1 3 0 {Rin}
* R2 1 3 {RFED}
.OP
* Analysis request
*2 .TF V(1) Vin
* 3-6 .TRAN {1/(freq*50)} {2/freq}
.AC DEC 20 1 1000MEG
* End the simulation
.END


