Simple RLC Circuit

* Circuit Description
* Low pass filter that passes the low freq and attenuate the high one
* Parameters

* Make avariable for cap and inductor
.PARAM C = 1p, L=1m

* Signal sources
* Add the voltage source between nodes 1 and 0(gnd)
* with AC mag=1 to make the gain=VOUT and phase=0
V1 1 0 AC 1
* Circuit elements
R1 1 2 100k
L1 2 3 1m
C1 3 0 1p
* Analysis request
* Run ac sweep from 1Hz to 100MEG with 10 pts per decade
.AC dec 10 1 100MEG
*** add line here ***
.PRINT AC V(1) V(3)
.PLOT AC V(1) V(3)

* Measure the peak
.MEAS AC PEAK max mag(V(3))

* Measure bandwidth using PEAK/sqrt(2)
.MEAS AC BW when mag(V(3))=PEAK/sqrt(2)

.End
